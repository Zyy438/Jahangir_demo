library verilog;
use verilog.vl_types.all;
entity soc_tb is
end soc_tb;
